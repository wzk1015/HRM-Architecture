`timescale 1ns / 1ps

module CPU(
		input [15:0] instr,
		input	[15:0] datain,
		input	[15:0] datain_final,
		input clk,
		input reset,
		output [15:0] pc,
		output [15:0] addr,
		output memWE
    );


endmodule
