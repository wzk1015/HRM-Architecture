`timescale 1ns / 1ps

module bridge(
    );


endmodule
