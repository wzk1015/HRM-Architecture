`timescale 1ns / 1ps

module inbox(
    );


endmodule
