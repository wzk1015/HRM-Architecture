`timescale 1ns / 1ps

module register(
		input [15:0] write_data,
		input clk,
		input reset,
		input WE,
		output [15:0] reg_data,
		output empty_reg
    );


endmodule
