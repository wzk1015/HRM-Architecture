`timescale 1ns / 1ps

module controller(
    );


endmodule
