`timescale 1ns / 1ps

module cp0(
    );


endmodule
