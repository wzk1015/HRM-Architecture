`timescale 1ns / 1ps

module npc(
		input [15:0] pc,
		input [15:0] cp0_pc,
		input [15:0] reg_val,
		input [11:0] j_addr,
		input [2:0] npc_sel,
		input exl,
		output [15:0] npc
    );


endmodule
